library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity HbbTV_Test_IP_v1_0 is
	generic (

		-- Parameters of Axi Slave Bus Interface S_AUDIO_AXIS
		C_S_AUDIO_AXIS_TDATA_WIDTH	: integer	:= 32;

		-- Parameters of Axi Master Bus Interface M_AUDIO_AXIS
		C_M_AUDIO_AXIS_TDATA_WIDTH	: integer	:= 32;

		-- Parameters of Axi Slave Bus Interface S_VIDEO_AXIS
		C_S_VIDEO_AXIS_TDATA_WIDTH	: integer	:= 32;

		-- Parameters of Axi Master Bus Interface M_VIDEO_AXIS
		C_M_VIDEO_AXIS_TDATA_WIDTH	: integer	:= 32;

		-- Parameters of Axi Slave Bus Interface S_CTRL_AXI
		C_S_CTRL_AXI_DATA_WIDTH	: integer	:= 32;
		C_S_CTRL_AXI_ADDR_WIDTH	: integer	:= 6
	);
	port (
		
		-- Ports of Axi Slave Bus Interface S_AUDIO_AXIS
		audio_aclk			: in std_logic;
		audio_aresetn		: in std_logic;
		s_audio_axis_tready	: out std_logic;
		s_audio_axis_tdata	: in std_logic_vector(C_S_AUDIO_AXIS_TDATA_WIDTH-1 downto 0);
		s_audio_axis_tlast	: in std_logic;
		s_audio_axis_tvalid	: in std_logic;

		-- Ports of Axi Master Bus Interface M_AUDIO_AXIS
		m_audio_axis_tvalid	: out std_logic;
		m_audio_axis_tdata	: out std_logic_vector(C_M_AUDIO_AXIS_TDATA_WIDTH-1 downto 0);
		m_audio_axis_tlast	: out std_logic;
		m_audio_axis_tready	: in std_logic;

		-- Ports of Axi Slave Bus Interface S_VIDEO_AXIS
		video_aclk			: in std_logic;
		video_aresetn		: in std_logic;
		s_video_axis_tready	: out std_logic;
		s_video_axis_tdata	: in std_logic_vector(C_S_VIDEO_AXIS_TDATA_WIDTH-1 downto 0);
		s_video_axis_tlast	: in std_logic;
		s_video_axis_tvalid	: in std_logic;
		s_video_axis_tuser	: in std_logic;

		-- Ports of Axi Master Bus Interface M_VIDEO_AXIS
		m_video_axis_tvalid	: out std_logic;
		m_video_axis_tdata	: out std_logic_vector(C_M_VIDEO_AXIS_TDATA_WIDTH-1 downto 0);
		m_video_axis_tlast	: out std_logic;
		m_video_axis_tuser	: out std_logic;
		m_video_axis_tready	: in std_logic;

		-- Ports of Axi Slave Bus Interface S_CTRL_AXI
		s_ctrl_axi_aclk	: in std_logic;
		s_ctrl_axi_aresetn	: in std_logic;
		s_ctrl_axi_awaddr	: in std_logic_vector(C_S_CTRL_AXI_ADDR_WIDTH-1 downto 0);
		s_ctrl_axi_awprot	: in std_logic_vector(2 downto 0);
		s_ctrl_axi_awvalid	: in std_logic;
		s_ctrl_axi_awready	: out std_logic;
		s_ctrl_axi_wdata	: in std_logic_vector(C_S_CTRL_AXI_DATA_WIDTH-1 downto 0);
		s_ctrl_axi_wstrb	: in std_logic_vector((C_S_CTRL_AXI_DATA_WIDTH/8)-1 downto 0);
		s_ctrl_axi_wvalid	: in std_logic;
		s_ctrl_axi_wready	: out std_logic;
		s_ctrl_axi_bresp	: out std_logic_vector(1 downto 0);
		s_ctrl_axi_bvalid	: out std_logic;
		s_ctrl_axi_bready	: in std_logic;
		s_ctrl_axi_araddr	: in std_logic_vector(C_S_CTRL_AXI_ADDR_WIDTH-1 downto 0);
		s_ctrl_axi_arprot	: in std_logic_vector(2 downto 0);
		s_ctrl_axi_arvalid	: in std_logic;
		s_ctrl_axi_arready	: out std_logic;
		s_ctrl_axi_rdata	: out std_logic_vector(C_S_CTRL_AXI_DATA_WIDTH-1 downto 0);
		s_ctrl_axi_rresp	: out std_logic_vector(1 downto 0);
		s_ctrl_axi_rvalid	: out std_logic;
		s_ctrl_axi_rready	: in std_logic
	);
end HbbTV_Test_IP_v1_0;

architecture arch_imp of HbbTV_Test_IP_v1_0 is

		signal HbbTV_audio_ready	: std_logic;
		signal HbbTV_video_ready	: std_logic;

		signal audio_data	: std_logic_vector(31 downto 0);
		signal audio_valid	: std_logic;
		signal audio_border	: std_logic_vector(31 downto 0);
		signal audio_ready	: std_logic;
		
		signal video_data	: std_logic_vector(31 downto 0);
		signal video_valid	: std_logic;
		signal video_last	: std_logic;
		signal video_sof	: std_logic;
		signal video_x1		: std_logic_vector(31 downto 0);
		signal video_x2		: std_logic_vector(31 downto 0);
		signal video_x3		: std_logic_vector(31 downto 0);
		signal video_x4		: std_logic_vector(31 downto 0);
		signal video_y1		: std_logic_vector(31 downto 0);
		signal video_y2		: std_logic_vector(31 downto 0);
		signal video_border	: std_logic_vector(31 downto 0);
		signal video_ready	: std_logic;
		
		signal synch_time	: std_logic_vector(15 downto 0);
	
	component HbbTV_Test is
		port	(
					iCLK					: in  std_logic;
					inRST					: in  std_logic;
					inPIXELS				: in  std_logic_vector(31 downto 0);
					inLAST_LINE				: in  std_logic;
					inVALID_PIXELS			: in  std_logic;
					inSTART_TRANSMISSION	: in  std_logic;
					inX1_COORDINATE			: in  std_logic_vector(31 downto 0);
					inX2_COORDINATE			: in  std_logic_vector(31 downto 0);
					inX3_COORDINATE			: in  std_logic_vector(31 downto 0);
					inX4_COORDINATE			: in  std_logic_vector(31 downto 0);
					inY1_COORDINATE			: in  std_logic_vector(31 downto 0);
					inY2_COORDINATE			: in  std_logic_vector(31 downto 0);
					inVIDEO_BORDER			: in  std_logic_vector(31 downto 0);
				
					inSAMPLES				: in  std_logic_vector(31 downto 0);
					inSAMPLES_VALID			: in  std_logic;
					inAUDIO_BORDER			: in  std_logic_vector(31 downto 0);
				
					outVIDEO_READY			: out std_logic;
					outAUDIO_READY			: out std_logic;
					outTIME					: out std_logic_vector(15 downto 0)	
				);
	end component HbbTV_Test;

	component HbbTV_Test_IP_v1_0_S_CTRL_AXI is
		generic (
		C_S_AXI_DATA_WIDTH	: integer	:= 32;
		C_S_AXI_ADDR_WIDTH	: integer	:= 6
		);
		port (
		
		outX1_COORDINATE	: out std_logic_vector(31 downto 0);
		outX2_COORDINATE	: out std_logic_vector(31 downto 0);
		outX3_COORDINATE	: out std_logic_vector(31 downto 0);
		outX4_COORDINATE	: out std_logic_vector(31 downto 0);
		outY1_COORDINATE	: out std_logic_vector(31 downto 0);
		outY2_COORDINATE	: out std_logic_vector(31 downto 0);
		outVIDEO_BORDER		: out std_logic_vector(31 downto 0);
		outAUDIO_BORDER		: out std_logic_vector(31 downto 0);
		inTIME				: in  std_logic_vector(15 downto 0);
		
		S_AXI_ACLK	: in std_logic;
		S_AXI_ARESETN	: in std_logic;
		S_AXI_AWADDR	: in std_logic_vector(C_S_AXI_ADDR_WIDTH-1 downto 0);
		S_AXI_AWPROT	: in std_logic_vector(2 downto 0);
		S_AXI_AWVALID	: in std_logic;
		S_AXI_AWREADY	: out std_logic;
		S_AXI_WDATA	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
		S_AXI_WSTRB	: in std_logic_vector((C_S_AXI_DATA_WIDTH/8)-1 downto 0);
		S_AXI_WVALID	: in std_logic;
		S_AXI_WREADY	: out std_logic;
		S_AXI_BRESP	: out std_logic_vector(1 downto 0);
		S_AXI_BVALID	: out std_logic;
		S_AXI_BREADY	: in std_logic;
		S_AXI_ARADDR	: in std_logic_vector(C_S_AXI_ADDR_WIDTH-1 downto 0);
		S_AXI_ARPROT	: in std_logic_vector(2 downto 0);
		S_AXI_ARVALID	: in std_logic;
		S_AXI_ARREADY	: out std_logic;
		S_AXI_RDATA	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
		S_AXI_RRESP	: out std_logic_vector(1 downto 0);
		S_AXI_RVALID	: out std_logic;
		S_AXI_RREADY	: in std_logic
		);
	end component HbbTV_Test_IP_v1_0_S_CTRL_AXI;

begin

-- Instantiation of Axi Bus Interface S_CTRL_AXI
HbbTV_Test_IP_v1_0_S_CTRL_AXI_inst : HbbTV_Test_IP_v1_0_S_CTRL_AXI
	generic map (
		C_S_AXI_DATA_WIDTH	=> C_S_CTRL_AXI_DATA_WIDTH,
		C_S_AXI_ADDR_WIDTH	=> C_S_CTRL_AXI_ADDR_WIDTH
	)
	port map (
		
		outX1_COORDINATE	=> video_x1,
		outX2_COORDINATE	=> video_x2,
		outX3_COORDINATE	=> video_x3,
		outX4_COORDINATE	=> video_x4,
		outY1_COORDINATE	=> video_y1,
		outY2_COORDINATE	=> video_y2,
		outVIDEO_BORDER		=> video_border,
		outAUDIO_BORDER		=> audio_border,
		inTIME				=> synch_time,
	
		S_AXI_ACLK	=> s_ctrl_axi_aclk,
		S_AXI_ARESETN	=> s_ctrl_axi_aresetn,
		S_AXI_AWADDR	=> s_ctrl_axi_awaddr,
		S_AXI_AWPROT	=> s_ctrl_axi_awprot,
		S_AXI_AWVALID	=> s_ctrl_axi_awvalid,
		S_AXI_AWREADY	=> s_ctrl_axi_awready,
		S_AXI_WDATA	=> s_ctrl_axi_wdata,
		S_AXI_WSTRB	=> s_ctrl_axi_wstrb,
		S_AXI_WVALID	=> s_ctrl_axi_wvalid,
		S_AXI_WREADY	=> s_ctrl_axi_wready,
		S_AXI_BRESP	=> s_ctrl_axi_bresp,
		S_AXI_BVALID	=> s_ctrl_axi_bvalid,
		S_AXI_BREADY	=> s_ctrl_axi_bready,
		S_AXI_ARADDR	=> s_ctrl_axi_araddr,
		S_AXI_ARPROT	=> s_ctrl_axi_arprot,
		S_AXI_ARVALID	=> s_ctrl_axi_arvalid,
		S_AXI_ARREADY	=> s_ctrl_axi_arready,
		S_AXI_RDATA	=> s_ctrl_axi_rdata,
		S_AXI_RRESP	=> s_ctrl_axi_rresp,
		S_AXI_RVALID	=> s_ctrl_axi_rvalid,
		S_AXI_RREADY	=> s_ctrl_axi_rready
	);

HbbTV_Test_inst:	HbbTV_Test port map	(
											iCLK					=> video_aclk,
											inRST					=> video_aresetn,
											inPIXELS				=> video_data,
											inLAST_LINE				=> video_last,
											inVALID_PIXELS			=> video_valid,
											inSTART_TRANSMISSION	=> video_sof,
											inX1_COORDINATE			=> video_x1,
											inX2_COORDINATE			=> video_x2,
											inX3_COORDINATE			=> video_x3,
											inX4_COORDINATE			=> video_x4,
											inY1_COORDINATE			=> video_y1,
											inY2_COORDINATE			=> video_y2,
											inVIDEO_BORDER			=> video_border,
											
											inSAMPLES				=> audio_data,
											inSAMPLES_VALID			=> audio_valid,
											inAUDIO_BORDER			=> audio_border,
											
											outVIDEO_READY			=> video_ready,
											outAUDIO_READY			=> audio_ready,
											outTIME					=> synch_time
										);
	audio_data	<= s_audio_axis_tdata;
	audio_valid	<= s_audio_axis_tvalid and m_audio_axis_tready;

	s_audio_axis_tready <= m_audio_axis_tready;

	m_audio_axis_tvalid <= s_audio_axis_tvalid;	
	m_audio_axis_tdata	<= audio_data;
	m_audio_axis_tlast	<= s_audio_axis_tlast;
	
	video_data	<= s_video_axis_tdata;
	video_valid	<= s_video_axis_tvalid and m_video_axis_tready;
	video_last	<= s_video_axis_tlast;
	video_sof	<= s_video_axis_tuser;
	
	s_video_axis_tready <= m_video_axis_tready;
	
	m_video_axis_tvalid	<= s_video_axis_tvalid;
	m_video_axis_tdata	<= video_data;
	m_video_axis_tlast	<= video_last;
	m_video_axis_tuser	<= video_sof;

end arch_imp;
